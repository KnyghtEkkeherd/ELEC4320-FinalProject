`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Name: Wiktor Kowalczyk
// Student ID: 20814029
// Email: wmkowalczyk@connect.ust.hk
//////////////////////////////////////////////////////////////////////////////////

module multiplier (
    input [31:0] A,
    input [31:0] B,
    input clk,
    output [63:0] P
);

    reg P;
    always @(posedge clk) begin

    end

endmodule
